// version_num
// this module contains the version number only
// format: 32'hYYMMDDHH
// Y  = Year  ('17' = 2017, '18' = 2018, '19' = 2019, '20' = 2020, , '21' = 2021, ...)
// M  = Month ('01..12' = Jan..Dec)
// DD = Day   (e.g. '01' = 01, '27' = 27, ...)
// DD = Hours (e.g. '01' = 01, '17' = 17, ...'23' = 23)
// Example: '17101209' = "2017 Oct. 12, 09 AM"
// Author: Dim Su
// Date: 20171012
// Do Not edit this file, its content to be changed automatically by appropriated TCL script

module version_num ( output [31:0] VERSION );
//VERSION:
assign VERSION = 32'h23062616;

endmodule






































































































































































































































































































































































































































































