`ifndef _define_led_driver_
`define _define_led_driver_

/******************************************************************************/
`define LED_DRIVER_MBI5153
//`define LED_DRIVER_MBI5124

/******************************************************************************/

`endif